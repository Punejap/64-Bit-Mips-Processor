
module top(
    input clk, reset;
);
